
module Pair(

    );
endmodule
